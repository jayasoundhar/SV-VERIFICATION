interface int_f();
  logic rst,clk;
  logic en;
  logic [3:0] data_in,data_out;
  logic full,empty;
endinterface
