interface int_f();
  logic [3:0]a;
  logic [3:0]b;
  logic cin;
  logic [3:0]sum;
  logic carry;
  
endinterface
