interface int_f();
  logic rst,clk;
  logic en;
  logic [7:0] data_in,data_out;
  logic [3:0] addr;
endinterface
