interface int_f();
  logic rst,clk;
  logic d;
  logic q,qb;
endinterface
