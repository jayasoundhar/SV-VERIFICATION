interface int_f();
  logic [3:0] out;
  logic rst,clk,s;
endinterface
